module Hex_PE_Cluster_quad(
    input  wire        clk,
    input  wire        reset_n,
    // 3 cặp IFM và Weightt
    input  wire [127:0]  Weight_0,
    input  wire [127:0]  Weight_1,
    input  wire [127:0]  Weight_2,
    input  wire [127:0]  Weight_3,
    input  wire [127:0]  IFM,
    // Tín hiệu điều khiển
    input  wire  [3:0] PE_reset,      
    input  wire  [3:0] PE_finish, 
    // Output
    output wire [7:0]  OFM_0,
    output wire [7:0]  OFM_1,
    output wire [7:0]  OFM_2,
    output wire [7:0]  OFM_3,
    output wire  [15:0]      valid
);
    Hex_PE instant_0 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),

        .Weight1 (Weight_0[7:0]),
        .Weight2 (Weight_0[15:8]),
        .Weight3 (Weight_0[23:16]),
        .Weight4 (Weight_0[31:24]),
        .Weight5 (Weight_0[39:32]),
        .Weight6 (Weight_0[47:40]),
        .Weight7 (Weight_0[55:48]),
        .Weight8 (Weight_0[63:56]),
        .Weight9 (Weight_0[71:64]),
        .Weight10(Weight_0[79:72]),
        .Weight11(Weight_0[87:80]),
        .Weight12(Weight_0[95:88]),
        .Weight13(Weight_0[103:96]),
        .Weight14(Weight_0[111:104]),
        .Weight15(Weight_0[119:112]),
        .Weight16(Weight_0[127:120]),

        .PE_reset(PE_reset[0]),
        .PE_finish(PE_finish[0]),
        .valid(valid[0]),
        .OFM(OFM_0)
    );
        Hex_PE instant_1 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),

        .Weight1 (Weight_1[7:0]),
        .Weight2 (Weight_1[15:8]),
        .Weight3 (Weight_1[23:16]),
        .Weight4 (Weight_1[31:24]),
        .Weight5 (Weight_1[39:32]),
        .Weight6 (Weight_1[47:40]),
        .Weight7 (Weight_1[55:48]),
        .Weight8 (Weight_1[63:56]),
        .Weight9 (Weight_1[71:64]),
        .Weight10(Weight_1[79:72]),
        .Weight11(Weight_1[87:80]),
        .Weight12(Weight_1[95:88]),
        .Weight13(Weight_1[103:96]),
        .Weight14(Weight_1[111:104]),
        .Weight15(Weight_1[119:112]),
        .Weight16(Weight_1[127:120]),

        .PE_reset(PE_reset[1]),
        .PE_finish(PE_finish[1]),
        .valid(valid[1]),
        .OFM(OFM_1)
    );
        Hex_PE instant_2 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),

        .Weight1 (Weight_2[7:0]),
        .Weight2 (Weight_2[15:8]),
        .Weight3 (Weight_2[23:16]),
        .Weight4 (Weight_2[31:24]),
        .Weight5 (Weight_2[39:32]),
        .Weight6 (Weight_2[47:40]),
        .Weight7 (Weight_2[55:48]),
        .Weight8 (Weight_2[63:56]),
        .Weight9 (Weight_2[71:64]),
        .Weight10(Weight_2[79:72]),
        .Weight11(Weight_2[87:80]),
        .Weight12(Weight_2[95:88]),
        .Weight13(Weight_2[103:96]),
        .Weight14(Weight_2[111:104]),
        .Weight15(Weight_2[119:112]),
        .Weight16(Weight_2[127:120]),

        .PE_reset(PE_reset[2]),
        .PE_finish(PE_finish[2]),
        .valid(valid[2]),
        .OFM(OFM_2)
    );
        Hex_PE instant_3 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),

        .Weight1 (Weight_3[7:0]),
        .Weight2 (Weight_3[15:8]),
        .Weight3 (Weight_3[23:16]),
        .Weight4 (Weight_3[31:24]),
        .Weight5 (Weight_3[39:32]),
        .Weight6 (Weight_3[47:40]),
        .Weight7 (Weight_3[55:48]),
        .Weight8 (Weight_3[63:56]),
        .Weight9 (Weight_3[71:64]),
        .Weight10(Weight_3[79:72]),
        .Weight11(Weight_3[87:80]),
        .Weight12(Weight_3[95:88]),
        .Weight13(Weight_3[103:96]),
        .Weight14(Weight_3[111:104]),
        .Weight15(Weight_3[119:112]),
        .Weight16(Weight_3[127:120]),
        .PE_reset(PE_reset[3]),
        .PE_finish(PE_finish[3]),
        .valid(valid[3]),
        .OFM(OFM_3)
    );
       
endmodule
module BRAM_General_weight #(
    parameter DATA_WIDTH_OUT    = 32,     // Số bit mỗi ô
    parameter DATA_WIDTH_IN    = 32,     // Số bit mỗi ô
    parameter DEPTH         = 8192,   // Tổng số ô nhớ
    parameter off_set_shift = 2       // Số bit dịch để truy cập theo word
)(
    input wire clk,
    input wire wr_rd_en,                               // Write enable
    input wire [$clog2(DEPTH)-1:0] wr_addr,            // Địa chỉ ghi
    input wire [$clog2(DEPTH*2**off_set_shift)-1:0] rd_addr,  // Địa chỉ đọc (địa chỉ byte → cần dịch)
    input wire [DATA_WIDTH_IN-1:0] data_in,               // Dữ liệu vào
    output reg [DATA_WIDTH_OUT-1:0] data_out               // Dữ liệu ra
    
);
    reg [127:0] data_load;
    // Khai báo RAM theo DEPTH
    (* ram_style = "block" *) reg [DATA_WIDTH_IN-1:0] bram [0:DEPTH-1];

    always @(posedge clk) begin
        if (wr_rd_en) begin
            bram[wr_addr] <= data_in;
        end
        
        case(rd_addr[3:2])
            2'b00: data_out <= bram[rd_addr >> off_set_shift] [31:0];
            2'b01: data_out <= bram[rd_addr >> off_set_shift] [63:32] ;
            2'b10: data_out <= bram[rd_addr >> off_set_shift] [95:64] ;
            2'b11: data_out <= bram[rd_addr >> off_set_shift] [127:96] ;
        endcase
    end
    // always_comb begin
    //     case(rd_addr[3:2])
    //         2'b00: data_out = data_load[31:0] ;
    //         2'b01: data_out = data_load[63:32] ;
    //         2'b10: data_out = data_load[95:64] ;
    //         2'b11: data_out = data_load[127:96] ;
    //     endcase
    // end
endmodule

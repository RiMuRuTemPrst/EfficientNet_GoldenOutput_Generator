module Hex_PE_cluster(
    input  wire        clk,
    input  wire        reset_n,
    // 3 cặp IFM và Weightt
    input  wire [127:0]  Weight_0,
    input  wire [127:0]  Weight_1,
    input  wire [127:0]  Weight_2,
    input  wire [127:0]  Weight_3,
    input  wire [127:0]  Weight_4,
    input  wire [127:0]  Weight_5,
    input  wire [127:0]  Weight_6,
    input  wire [127:0]  Weight_7,
    input  wire [127:0]  Weight_8,
    input  wire [127:0]  Weight_9,
    input  wire [127:0]  Weight_10,
    input  wire [127:0]  Weight_11,
    input  wire [127:0]  Weight_12,
    input  wire [127:0]  Weight_13,
    input  wire [127:0]  Weight_14,
    input  wire [127:0]  Weight_15,
    input  wire [127:0]  IFM,
    // Tín hiệu điều khiển
    input  wire  [15:0] PE_reset,      
    input  wire  [15:0] PE_finish, 
    // Output
    output wire [7:0]  OFM_0,
    output wire [7:0]  OFM_1,
    output wire [7:0]  OFM_2,
    output wire [7:0]  OFM_3,
    output wire [7:0]  OFM_4,
    output wire [7:0]  OFM_5,
    output wire [7:0]  OFM_6,
    output wire [7:0]  OFM_7,
    output wire [7:0]  OFM_8,
    output wire [7:0]  OFM_9,
    output wire [7:0]  OFM_10,
    output wire [7:0]  OFM_11,
    output wire [7:0]  OFM_12,
    output wire [7:0]  OFM_13,
    output wire [7:0]  OFM_14,
    output wire [7:0]  OFM_15,
    output wire [7:0]  OFM_16,
    output wire  [15:0]      valid
);
    Hex_PE instant_0 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_0[7:0]),
        .Weight2 (Weight_0[15:8]),
        .Weight3 (Weight_0[23:16]),
        .Weight4 (Weight_0[31:24]),
        .Weight5 (Weight_0[39:32]),
        .Weight6 (Weight_0[47:40]),
        .Weight7 (Weight_0[55:48]),
        .Weight8 (Weight_0[63:56]),
        .Weight9 (Weight_0[71:64]),
        .Weight10(Weight_0[79:72]),
        .Weight11(Weight_0[87:80]),
        .Weight12(Weight_0[95:88]),
        .Weight13(Weight_0[103:96]),
        .Weight14(Weight_0[111:104]),
        .Weight15(Weight_0[119:112]),
        .Weight16(Weight_0[127:120]),
        .PE_reset(PE_reset[0]),
        .PE_finish(PE_finish[0]),
        .valid(valid[0]),
        .OFM(OFM_0)
    );
        Hex_PE instant_1 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_1[7:0]),
        .Weight2 (Weight_1[15:8]),
        .Weight3 (Weight_1[23:16]),
        .Weight4 (Weight_1[31:24]),
        .Weight5 (Weight_1[39:32]),
        .Weight6 (Weight_1[47:40]),
        .Weight7 (Weight_1[55:48]),
        .Weight8 (Weight_1[63:56]),
        .Weight9 (Weight_1[71:64]),
        .Weight10(Weight_1[79:72]),
        .Weight11(Weight_1[87:80]),
        .Weight12(Weight_1[95:88]),
        .Weight13(Weight_1[103:96]),
        .Weight14(Weight_1[111:104]),
        .Weight15(Weight_1[119:112]),
        .Weight16(Weight_1[127:120]),
        .PE_reset(PE_reset[1]),
        .PE_finish(PE_finish[1]),
        .valid(valid[1]),
        .OFM(OFM_1)
    );
        Hex_PE instant_2 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_2[7:0]),
        .Weight2 (Weight_2[15:8]),
        .Weight3 (Weight_2[23:16]),
        .Weight4 (Weight_2[31:24]),
        .Weight5 (Weight_2[39:32]),
        .Weight6 (Weight_2[47:40]),
        .Weight7 (Weight_2[55:48]),
        .Weight8 (Weight_2[63:56]),
        .Weight9 (Weight_2[71:64]),
        .Weight10(Weight_2[79:72]),
        .Weight11(Weight_2[87:80]),
        .Weight12(Weight_2[95:88]),
        .Weight13(Weight_2[103:96]),
        .Weight14(Weight_2[111:104]),
        .Weight15(Weight_2[119:112]),
        .Weight16(Weight_2[127:120]),
        .PE_reset(PE_reset[2]),
        .PE_finish(PE_finish[2]),
        .valid(valid[2]),
        .OFM(OFM_2)
    );
        Hex_PE instant_3 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_3[7:0]),
        .Weight2 (Weight_3[15:8]),
        .Weight3 (Weight_3[23:16]),
        .Weight4 (Weight_3[31:24]),
        .Weight5 (Weight_3[39:32]),
        .Weight6 (Weight_3[47:40]),
        .Weight7 (Weight_3[55:48]),
        .Weight8 (Weight_3[63:56]),
        .Weight9 (Weight_3[71:64]),
        .Weight10(Weight_3[79:72]),
        .Weight11(Weight_3[87:80]),
        .Weight12(Weight_3[95:88]),
        .Weight13(Weight_3[103:96]),
        .Weight14(Weight_3[111:104]),
        .Weight15(Weight_3[119:112]),
        .Weight16(Weight_3[127:120]),
        .PE_reset(PE_reset[3]),
        .PE_finish(PE_finish[3]),
        .valid(valid[3]),
        .OFM(OFM_3)
    );
        Hex_PE instant_4 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_4[7:0]),
        .Weight2 (Weight_4[15:8]),
        .Weight3 (Weight_4[23:16]),
        .Weight4 (Weight_4[31:24]),
        .Weight5 (Weight_4[39:32]),
        .Weight6 (Weight_4[47:40]),
        .Weight7 (Weight_4[55:48]),
        .Weight8 (Weight_4[63:56]),
        .Weight9 (Weight_4[71:64]),
        .Weight10(Weight_4[79:72]),
        .Weight11(Weight_4[87:80]),
        .Weight12(Weight_4[95:88]),
        .Weight13(Weight_4[103:96]),
        .Weight14(Weight_4[111:104]),
        .Weight15(Weight_4[119:112]),
        .Weight16(Weight_4[127:120]),
        .PE_reset(PE_reset[4]),
        .PE_finish(PE_finish[4]),
        .valid(valid[4]),
        .OFM(OFM_4)
    );
        Hex_PE instant_5 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_5[7:0]),
        .Weight2 (Weight_5[15:8]),
        .Weight3 (Weight_5[23:16]),
        .Weight4 (Weight_5[31:24]),
        .Weight5 (Weight_5[39:32]),
        .Weight6 (Weight_5[47:40]),
        .Weight7 (Weight_5[55:48]),
        .Weight8 (Weight_5[63:56]),
        .Weight9 (Weight_5[71:64]),
        .Weight10(Weight_5[79:72]),
        .Weight11(Weight_5[87:80]),
        .Weight12(Weight_5[95:88]),
        .Weight13(Weight_5[103:96]),
        .Weight14(Weight_5[111:104]),
        .Weight15(Weight_5[119:112]),
        .Weight16(Weight_5[127:120]),
        .PE_reset(PE_reset[5]),
        .PE_finish(PE_finish[5]),
        .valid(valid[5]),
        .OFM(OFM_5)
    );
        Hex_PE instant_6 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_6[7:0]),
        .Weight2 (Weight_6[15:8]),
        .Weight3 (Weight_6[23:16]),
        .Weight4 (Weight_6[31:24]),
        .Weight5 (Weight_6[39:32]),
        .Weight6 (Weight_6[47:40]),
        .Weight7 (Weight_6[55:48]),
        .Weight8 (Weight_6[63:56]),
        .Weight9 (Weight_6[71:64]),
        .Weight10(Weight_6[79:72]),
        .Weight11(Weight_6[87:80]),
        .Weight12(Weight_6[95:88]),
        .Weight13(Weight_6[103:96]),
        .Weight14(Weight_6[111:104]),
        .Weight15(Weight_6[119:112]),
        .Weight16(Weight_6[127:120]),
        .PE_reset(PE_reset[6]),
        .PE_finish(PE_finish[6]),
        .valid(valid[6]),
        .OFM(OFM_6)
    );
        Hex_PE instant_7 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_7[7:0]),
        .Weight2 (Weight_7[15:8]),
        .Weight3 (Weight_7[23:16]),
        .Weight4 (Weight_7[31:24]),
        .Weight5 (Weight_7[39:32]),
        .Weight6 (Weight_7[47:40]),
        .Weight7 (Weight_7[55:48]),
        .Weight8 (Weight_7[63:56]),
        .Weight9 (Weight_7[71:64]),
        .Weight10(Weight_7[79:72]),
        .Weight11(Weight_7[87:80]),
        .Weight12(Weight_7[95:88]),
        .Weight13(Weight_7[103:96]),
        .Weight14(Weight_7[111:104]),
        .Weight15(Weight_7[119:112]),
        .Weight16(Weight_7[127:120]),
        .PE_reset(PE_reset[7]),
        .PE_finish(PE_finish[7]),
        .valid(valid[7]),
        .OFM(OFM_7)
    );
        Hex_PE instant_8 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_8[7:0]),
        .Weight2 (Weight_8[15:8]),
        .Weight3 (Weight_8[23:16]),
        .Weight4 (Weight_8[31:24]),
        .Weight5 (Weight_8[39:32]),
        .Weight6 (Weight_8[47:40]),
        .Weight7 (Weight_8[55:48]),
        .Weight8 (Weight_8[63:56]),
        .Weight9 (Weight_8[71:64]),
        .Weight10(Weight_8[79:72]),
        .Weight11(Weight_8[87:80]),
        .Weight12(Weight_8[95:88]),
        .Weight13(Weight_8[103:96]),
        .Weight14(Weight_8[111:104]),
        .Weight15(Weight_8[119:112]),
        .Weight16(Weight_8[127:120]),
        .PE_reset(PE_reset[8]),
        .PE_finish(PE_finish[8]),
        .valid(valid[8]),
        .OFM(OFM_8)
    );
        Hex_PE instant_9 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_9[7:0]),
        .Weight2 (Weight_9[15:8]),
        .Weight3 (Weight_9[23:16]),
        .Weight4 (Weight_9[31:24]),
        .Weight5 (Weight_9[39:32]),
        .Weight6 (Weight_9[47:40]),
        .Weight7 (Weight_9[55:48]),
        .Weight8 (Weight_9[63:56]),
        .Weight9 (Weight_9[71:64]),
        .Weight10(Weight_9[79:72]),
        .Weight11(Weight_9[87:80]),
        .Weight12(Weight_9[95:88]),
        .Weight13(Weight_9[103:96]),
        .Weight14(Weight_9[111:104]),
        .Weight15(Weight_9[119:112]),
        .Weight16(Weight_9[127:120]),
        .PE_reset(PE_reset[9]),
        .PE_finish(PE_finish[9]),
        .valid(valid[9]),
        .OFM(OFM_9)
    );
        Hex_PE instant_10 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_10[7:0]),
        .Weight2 (Weight_10[15:8]),
        .Weight3 (Weight_10[23:16]),
        .Weight4 (Weight_10[31:24]),
        .Weight5 (Weight_10[39:32]),
        .Weight6 (Weight_10[47:40]),
        .Weight7 (Weight_10[55:48]),
        .Weight8 (Weight_10[63:56]),
        .Weight9 (Weight_10[71:64]),
        .Weight10(Weight_10[79:72]),
        .Weight11(Weight_10[87:80]),
        .Weight12(Weight_10[95:88]),
        .Weight13(Weight_10[103:96]),
        .Weight14(Weight_10[111:104]),
        .Weight15(Weight_10[119:112]),
        .Weight16(Weight_10[127:120]),
        .PE_reset(PE_reset[10]),
        .PE_finish(PE_finish[10]),
        .valid(valid[10]),
        .OFM(OFM_10)
    );
        Hex_PE instant_11 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_11[7:0]),
        .Weight2 (Weight_11[15:8]),
        .Weight3 (Weight_11[23:16]),
        .Weight4 (Weight_11[31:24]),
        .Weight5 (Weight_11[39:32]),
        .Weight6 (Weight_11[47:40]),
        .Weight7 (Weight_11[55:48]),
        .Weight8 (Weight_11[63:56]),
        .Weight9 (Weight_11[71:64]),
        .Weight10(Weight_11[79:72]),
        .Weight11(Weight_11[87:80]),
        .Weight12(Weight_11[95:88]),
        .Weight13(Weight_11[103:96]),
        .Weight14(Weight_11[111:104]),
        .Weight15(Weight_11[119:112]),
        .Weight16(Weight_11[127:120]),
        .PE_reset(PE_reset[11]),
        .PE_finish(PE_finish[11]),
        .valid(valid[11]),
        .OFM(OFM_11)
    );
        Hex_PE instant_12 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_12[7:0]),
        .Weight2 (Weight_12[15:8]),
        .Weight3 (Weight_12[23:16]),
        .Weight4 (Weight_12[31:24]),
        .Weight5 (Weight_12[39:32]),
        .Weight6 (Weight_12[47:40]),
        .Weight7 (Weight_12[55:48]),
        .Weight8 (Weight_12[63:56]),
        .Weight9 (Weight_12[71:64]),
        .Weight10(Weight_12[79:72]),
        .Weight11(Weight_12[87:80]),
        .Weight12(Weight_12[95:88]),
        .Weight13(Weight_12[103:96]),
        .Weight14(Weight_12[111:104]),
        .Weight15(Weight_12[119:112]),
        .Weight16(Weight_12[127:120]),
        .PE_reset(PE_reset[12]),
        .PE_finish(PE_finish[12]),
        .valid(valid[12]),
        .OFM(OFM_12)
    );
           Hex_PE instant_13 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_13[7:0]),
        .Weight2 (Weight_13[15:8]),
        .Weight3 (Weight_13[23:16]),
        .Weight4 (Weight_13[31:24]),
        .Weight5 (Weight_13[39:32]),
        .Weight6 (Weight_13[47:40]),
        .Weight7 (Weight_13[55:48]),
        .Weight8 (Weight_13[63:56]),
        .Weight9 (Weight_13[71:64]),
        .Weight10(Weight_13[79:72]),
        .Weight11(Weight_13[87:80]),
        .Weight12(Weight_13[95:88]),
        .Weight13(Weight_13[103:96]),
        .Weight14(Weight_13[111:104]),
        .Weight15(Weight_13[119:112]),
        .Weight16(Weight_13[127:120]),
        .PE_reset(PE_reset[13]),
        .PE_finish(PE_finish[13]),
        .valid(valid[13]),
        .OFM(OFM_13)
    );
            Hex_PE instant_14 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_14[7:0]),
        .Weight2 (Weight_14[15:8]),
        .Weight3 (Weight_14[23:16]),
        .Weight4 (Weight_14[31:24]),
        .Weight5 (Weight_14[39:32]),
        .Weight6 (Weight_14[47:40]),
        .Weight7 (Weight_14[55:48]),
        .Weight8 (Weight_14[63:56]),
        .Weight9 (Weight_14[71:64]),
        .Weight10(Weight_14[79:72]),
        .Weight11(Weight_14[87:80]),
        .Weight12(Weight_14[95:88]),
        .Weight13(Weight_14[103:96]),
        .Weight14(Weight_14[111:104]),
        .Weight15(Weight_14[119:112]),
        .Weight16(Weight_14[127:120]),
        .PE_reset(PE_reset[14]),
        .PE_finish(PE_finish[14]),
        .valid(valid[14]),
        .OFM(OFM_14)
    );
            Hex_PE instant_15 (
        .clk(clk),
        .reset_n(reset_n),
        .IFM1 (IFM[7:0]),
        .IFM2 (IFM[15:8]),
        .IFM3 (IFM[23:16]),
        .IFM4 (IFM[31:24]),
        .IFM5 (IFM[39:32]),
        .IFM6 (IFM[47:40]),
        .IFM7 (IFM[55:48]),
        .IFM8 (IFM[63:56]),
        .IFM9 (IFM[71:64]),
        .IFM10(IFM[79:72]),
        .IFM11(IFM[87:80]),
        .IFM12(IFM[95:88]),
        .IFM13(IFM[103:96]),
        .IFM14(IFM[111:104]),
        .IFM15(IFM[119:112]),
        .IFM16(IFM[127:120]),
        .Weight1 (Weight_15[7:0]),
        .Weight2 (Weight_15[15:8]),
        .Weight3 (Weight_15[23:16]),
        .Weight4 (Weight_15[31:24]),
        .Weight5 (Weight_15[39:32]),
        .Weight6 (Weight_15[47:40]),
        .Weight7 (Weight_15[55:48]),
        .Weight8 (Weight_15[63:56]),
        .Weight9 (Weight_15[71:64]),
        .Weight10(Weight_15[79:72]),
        .Weight11(Weight_15[87:80]),
        .Weight12(Weight_15[95:88]),
        .Weight13(Weight_15[103:96]),
        .Weight14(Weight_15[111:104]),
        .Weight15(Weight_15[119:112]),
        .Weight16(Weight_15[127:120]),
        .PE_reset(PE_reset[15]),
        .PE_finish(PE_finish[15]),
        .valid(valid[15]),
        .OFM(OFM_15)
    );

endmodule